module verifica_len_out(
  input logic [2:0] len_out,
  output logic ack_in 
);

  
