module verifica_len_out(
  input logic []len_out,
  output logic ack_in 
);

  
