module fila(
    input [7:0] data_in,
    input enqueue_in,
    input dequeue_in
    
    input reset,
    input clock,
    
    output data_out,
    output len_out,
);
